* NGSPICE file created from cs.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_WUV6BX a_26_n438# a_207_n350# a_n29_n350# a_89_n350#
+ a_n210_n438# a_n564_n438# a_n721_n524# a_n92_n438# a_n501_n350# a_380_n438# a_n446_n438#
+ a_561_n350# a_n383_n350# a_262_n438# a_n328_n438# a_443_n350# a_n265_n350# a_n619_n350#
+ a_498_n438# a_144_n438# a_325_n350# a_n147_n350#
X0 a_325_n350# a_262_n438# a_207_n350# a_n721_n524# sky130_fd_pr__nfet_01v8 ad=0.507 pd=3.79 as=0.507 ps=3.79 w=3.5 l=0.3
X1 a_n265_n350# a_n328_n438# a_n383_n350# a_n721_n524# sky130_fd_pr__nfet_01v8 ad=0.507 pd=3.79 as=0.507 ps=3.79 w=3.5 l=0.3
X2 a_561_n350# a_498_n438# a_443_n350# a_n721_n524# sky130_fd_pr__nfet_01v8 ad=1.01 pd=7.58 as=0.507 ps=3.79 w=3.5 l=0.3
X3 a_89_n350# a_26_n438# a_n29_n350# a_n721_n524# sky130_fd_pr__nfet_01v8 ad=0.507 pd=3.79 as=0.507 ps=3.79 w=3.5 l=0.3
X4 a_207_n350# a_144_n438# a_89_n350# a_n721_n524# sky130_fd_pr__nfet_01v8 ad=0.507 pd=3.79 as=0.507 ps=3.79 w=3.5 l=0.3
X5 a_n501_n350# a_n564_n438# a_n619_n350# a_n721_n524# sky130_fd_pr__nfet_01v8 ad=0.507 pd=3.79 as=1.01 ps=7.58 w=3.5 l=0.3
X6 a_n147_n350# a_n210_n438# a_n265_n350# a_n721_n524# sky130_fd_pr__nfet_01v8 ad=0.507 pd=3.79 as=0.507 ps=3.79 w=3.5 l=0.3
X7 a_443_n350# a_380_n438# a_325_n350# a_n721_n524# sky130_fd_pr__nfet_01v8 ad=0.507 pd=3.79 as=0.507 ps=3.79 w=3.5 l=0.3
X8 a_n383_n350# a_n446_n438# a_n501_n350# a_n721_n524# sky130_fd_pr__nfet_01v8 ad=0.507 pd=3.79 as=0.507 ps=3.79 w=3.5 l=0.3
X9 a_n29_n350# a_n92_n438# a_n147_n350# a_n721_n524# sky130_fd_pr__nfet_01v8 ad=0.507 pd=3.79 as=0.507 ps=3.79 w=3.5 l=0.3
C0 a_26_n438# a_144_n438# 0.112f
C1 a_n29_n350# a_89_n350# 0.418f
C2 a_26_n438# a_n92_n438# 0.112f
C3 a_561_n350# a_443_n350# 0.418f
C4 a_89_n350# a_207_n350# 0.418f
C5 a_561_n350# a_498_n438# 0.0308f
C6 a_n147_n350# a_n210_n438# 0.0308f
C7 a_n29_n350# a_n92_n438# 0.0308f
C8 a_207_n350# a_144_n438# 0.0308f
C9 a_n265_n350# a_n383_n350# 0.418f
C10 a_n501_n350# a_n383_n350# 0.418f
C11 a_n501_n350# a_n564_n438# 0.0308f
C12 a_443_n350# a_498_n438# 0.0308f
C13 a_n265_n350# a_n147_n350# 0.418f
C14 a_n446_n438# a_n328_n438# 0.112f
C15 a_n265_n350# a_n210_n438# 0.0308f
C16 a_262_n438# a_144_n438# 0.112f
C17 a_380_n438# a_325_n350# 0.0308f
C18 a_n29_n350# a_26_n438# 0.0308f
C19 a_n147_n350# a_n92_n438# 0.0308f
C20 a_325_n350# a_207_n350# 0.418f
C21 a_n210_n438# a_n92_n438# 0.112f
C22 a_n383_n350# a_n446_n438# 0.0308f
C23 a_n446_n438# a_n564_n438# 0.112f
C24 a_n564_n438# a_n619_n350# 0.0308f
C25 a_262_n438# a_325_n350# 0.0308f
C26 a_380_n438# a_262_n438# 0.112f
C27 a_89_n350# a_144_n438# 0.0308f
C28 a_n383_n350# a_n328_n438# 0.0308f
C29 a_262_n438# a_207_n350# 0.0308f
C30 a_325_n350# a_443_n350# 0.418f
C31 a_380_n438# a_443_n350# 0.0308f
C32 a_n29_n350# a_n147_n350# 0.418f
C33 a_n210_n438# a_n328_n438# 0.112f
C34 a_n501_n350# a_n446_n438# 0.0308f
C35 a_n501_n350# a_n619_n350# 0.418f
C36 a_380_n438# a_498_n438# 0.112f
C37 a_89_n350# a_26_n438# 0.0308f
C38 a_n265_n350# a_n328_n438# 0.0308f
C39 a_561_n350# a_n721_n524# 0.398f
C40 a_443_n350# a_n721_n524# 0.0725f
C41 a_325_n350# a_n721_n524# 0.0725f
C42 a_207_n350# a_n721_n524# 0.0725f
C43 a_89_n350# a_n721_n524# 0.0725f
C44 a_n29_n350# a_n721_n524# 0.0725f
C45 a_n147_n350# a_n721_n524# 0.0725f
C46 a_n265_n350# a_n721_n524# 0.0725f
C47 a_n383_n350# a_n721_n524# 0.0725f
C48 a_n501_n350# a_n721_n524# 0.0725f
C49 a_n619_n350# a_n721_n524# 0.398f
C50 a_498_n438# a_n721_n524# 0.285f
C51 a_380_n438# a_n721_n524# 0.218f
C52 a_262_n438# a_n721_n524# 0.218f
C53 a_144_n438# a_n721_n524# 0.218f
C54 a_26_n438# a_n721_n524# 0.218f
C55 a_n92_n438# a_n721_n524# 0.218f
C56 a_n210_n438# a_n721_n524# 0.218f
C57 a_n328_n438# a_n721_n524# 0.218f
C58 a_n446_n438# a_n721_n524# 0.218f
C59 a_n564_n438# a_n721_n524# 0.285f
.ends

.subckt sky130_fd_pr__res_xhigh_po_2p85_RYTYPJ a_n285_n575# a_n415_n705# a_n285_143#
X0 a_n285_143# a_n285_n575# a_n415_n705# sky130_fd_pr__res_xhigh_po_2p85 l=1.43
C0 a_n285_143# a_n285_n575# 0.117f
C1 a_n285_n575# a_n415_n705# 1.05f
C2 a_n285_143# a_n415_n705# 1.05f
.ends

.subckt cs inp out vdd vss
XXM1 inp vss vss out inp inp vss inp vss inp inp out out inp inp vss vss out inp inp
+ out out sky130_fd_pr__nfet_01v8_WUV6BX
Xsky130_fd_pr__res_xhigh_po_2p85_RYTYPJ_0 out vss vdd sky130_fd_pr__res_xhigh_po_2p85_RYTYPJ
C0 inp vdd 6.45e-19
C1 vss vdd 0.0435f
C2 inp out 1.17f
C3 vss out 1.43f
C4 vss inp 1.21f
C5 out vdd 0.073f
C6 vss 0 0.935f
C7 vdd 0 1.75f
C8 out 0 3.1f
C9 inp 0 2.94f
.ends

