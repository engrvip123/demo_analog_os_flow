* NGSPICE file created from cs.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_2p85_53STJD a_n285_n559# a_n415_n689# a_n285_127#
X0 a_n285_127# a_n285_n559# a_n415_n689# sky130_fd_pr__res_xhigh_po_2p85 l=1.43
C0 a_n285_n559# a_n285_127# 0.129933f
C1 a_n285_n559# a_n415_n689# 1.03823f
C2 a_n285_127# a_n415_n689# 1.03823f
.ends

.subckt sky130_fd_pr__nfet_01v8_WUV6BX a_26_n438# a_207_n350# a_n29_n350# a_89_n350#
+ a_n210_n438# a_n564_n438# a_n721_n524# a_n92_n438# a_n501_n350# a_380_n438# a_n446_n438#
+ a_561_n350# a_n383_n350# a_262_n438# a_n328_n438# a_443_n350# a_n265_n350# a_n619_n350#
+ a_498_n438# a_144_n438# a_325_n350# a_n147_n350#
X0 a_325_n350# a_262_n438# a_207_n350# a_n721_n524# sky130_fd_pr__nfet_01v8 ad=0.5075 pd=3.79 as=0.5075 ps=3.79 w=3.5 l=0.3
X1 a_n265_n350# a_n328_n438# a_n383_n350# a_n721_n524# sky130_fd_pr__nfet_01v8 ad=0.5075 pd=3.79 as=0.5075 ps=3.79 w=3.5 l=0.3
X2 a_561_n350# a_498_n438# a_443_n350# a_n721_n524# sky130_fd_pr__nfet_01v8 ad=1.015 pd=7.58 as=0.5075 ps=3.79 w=3.5 l=0.3
X3 a_89_n350# a_26_n438# a_n29_n350# a_n721_n524# sky130_fd_pr__nfet_01v8 ad=0.5075 pd=3.79 as=0.5075 ps=3.79 w=3.5 l=0.3
X4 a_207_n350# a_144_n438# a_89_n350# a_n721_n524# sky130_fd_pr__nfet_01v8 ad=0.5075 pd=3.79 as=0.5075 ps=3.79 w=3.5 l=0.3
X5 a_n501_n350# a_n564_n438# a_n619_n350# a_n721_n524# sky130_fd_pr__nfet_01v8 ad=0.5075 pd=3.79 as=1.015 ps=7.58 w=3.5 l=0.3
X6 a_n147_n350# a_n210_n438# a_n265_n350# a_n721_n524# sky130_fd_pr__nfet_01v8 ad=0.5075 pd=3.79 as=0.5075 ps=3.79 w=3.5 l=0.3
X7 a_443_n350# a_380_n438# a_325_n350# a_n721_n524# sky130_fd_pr__nfet_01v8 ad=0.5075 pd=3.79 as=0.5075 ps=3.79 w=3.5 l=0.3
X8 a_n383_n350# a_n446_n438# a_n501_n350# a_n721_n524# sky130_fd_pr__nfet_01v8 ad=0.5075 pd=3.79 as=0.5075 ps=3.79 w=3.5 l=0.3
X9 a_n29_n350# a_n92_n438# a_n147_n350# a_n721_n524# sky130_fd_pr__nfet_01v8 ad=0.5075 pd=3.79 as=0.5075 ps=3.79 w=3.5 l=0.3
C0 a_n210_n438# a_n265_n350# 0.030826f
C1 a_498_n438# a_380_n438# 0.112166f
C2 a_144_n438# a_262_n438# 0.112166f
C3 a_443_n350# a_380_n438# 0.030826f
C4 a_262_n438# a_380_n438# 0.112166f
C5 a_n265_n350# a_n147_n350# 0.417904f
C6 a_207_n350# a_89_n350# 0.417904f
C7 a_325_n350# a_207_n350# 0.417904f
C8 a_n446_n438# a_n564_n438# 0.112166f
C9 a_89_n350# a_26_n438# 0.030826f
C10 a_n210_n438# a_n92_n438# 0.112166f
C11 a_498_n438# a_561_n350# 0.030826f
C12 a_n446_n438# a_n501_n350# 0.030826f
C13 a_561_n350# a_443_n350# 0.417904f
C14 a_207_n350# a_144_n438# 0.030826f
C15 a_n564_n438# a_n501_n350# 0.030826f
C16 a_n92_n438# a_n147_n350# 0.030826f
C17 a_498_n438# a_443_n350# 0.030826f
C18 a_26_n438# a_n92_n438# 0.112166f
C19 a_26_n438# a_144_n438# 0.112166f
C20 a_n328_n438# a_n383_n350# 0.030826f
C21 a_89_n350# a_144_n438# 0.030826f
C22 a_325_n350# a_380_n438# 0.030826f
C23 a_n328_n438# a_n210_n438# 0.112166f
C24 a_n29_n350# a_n147_n350# 0.417904f
C25 a_207_n350# a_262_n438# 0.030826f
C26 a_26_n438# a_n29_n350# 0.030826f
C27 a_n619_n350# a_n564_n438# 0.030826f
C28 a_89_n350# a_n29_n350# 0.417904f
C29 a_n328_n438# a_n265_n350# 0.030826f
C30 a_n328_n438# a_n446_n438# 0.112166f
C31 a_n619_n350# a_n501_n350# 0.417904f
C32 a_n383_n350# a_n265_n350# 0.417904f
C33 a_n446_n438# a_n383_n350# 0.030826f
C34 a_325_n350# a_443_n350# 0.417904f
C35 a_325_n350# a_262_n438# 0.030826f
C36 a_n210_n438# a_n147_n350# 0.030826f
C37 a_n383_n350# a_n501_n350# 0.417904f
C38 a_n92_n438# a_n29_n350# 0.030826f
C39 a_561_n350# a_n721_n524# 0.397781f
C40 a_443_n350# a_n721_n524# 0.072511f
C41 a_325_n350# a_n721_n524# 0.072511f
C42 a_207_n350# a_n721_n524# 0.072511f
C43 a_89_n350# a_n721_n524# 0.072511f
C44 a_n29_n350# a_n721_n524# 0.072511f
C45 a_n147_n350# a_n721_n524# 0.072511f
C46 a_n265_n350# a_n721_n524# 0.072511f
C47 a_n383_n350# a_n721_n524# 0.072511f
C48 a_n501_n350# a_n721_n524# 0.072511f
C49 a_n619_n350# a_n721_n524# 0.397781f
C50 a_498_n438# a_n721_n524# 0.284614f
C51 a_380_n438# a_n721_n524# 0.218475f
C52 a_262_n438# a_n721_n524# 0.21835f
C53 a_144_n438# a_n721_n524# 0.218301f
C54 a_26_n438# a_n721_n524# 0.218283f
C55 a_n92_n438# a_n721_n524# 0.218283f
C56 a_n210_n438# a_n721_n524# 0.218301f
C57 a_n328_n438# a_n721_n524# 0.21835f
C58 a_n446_n438# a_n721_n524# 0.218475f
C59 a_n564_n438# a_n721_n524# 0.284614f
.ends

.subckt cs out inp vdd vss
XXR2 out vss vdd sky130_fd_pr__res_xhigh_po_2p85_53STJD
XXM1 inp vss vss out inp inp vss inp vss inp inp out out inp inp vss vss out inp inp
+ out out sky130_fd_pr__nfet_01v8_WUV6BX
C0 inp vdd 6.26e-19
C1 out vdd 0.078799f
C2 out inp 1.262959f
C3 inp vss 4.116509f
C4 out vss 5.397398f
C5 vdd vss 1.452687f
.ends

