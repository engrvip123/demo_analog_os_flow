magic
tech sky130A
magscale 1 2
timestamp 1705487333
<< pwell >>
rect 984 1420 1128 1482
<< locali >>
rect 350 1602 394 2044
<< viali >>
rect 426 552 1056 618
<< metal1 >>
rect 506 2786 988 3674
rect 506 2072 516 2444
rect 1022 2072 1032 2444
rect 1550 1686 1560 1976
rect 1870 1686 1880 1976
rect -158 1540 1182 1542
rect -158 1486 1276 1540
rect -158 1485 1182 1486
rect -153 1188 -95 1485
rect -300 988 -95 1188
rect 62 1136 72 1444
rect 142 1136 152 1444
rect 310 1136 320 1444
rect 390 1136 400 1444
rect 546 1136 556 1444
rect 626 1136 636 1444
rect 782 1136 792 1444
rect 862 1136 872 1444
rect 1016 1136 1026 1444
rect 1096 1136 1106 1444
rect 1254 1136 1264 1444
rect 1334 1136 1344 1444
rect -153 770 -95 988
rect -154 726 -94 770
rect 184 766 194 1042
rect 262 766 272 1042
rect 428 768 438 1044
rect 506 768 516 1044
rect 666 768 676 1044
rect 744 768 754 1044
rect 902 774 912 1050
rect 980 774 990 1050
rect 1136 770 1146 1046
rect 1214 770 1224 1046
rect -154 678 1280 726
rect 414 618 1068 624
rect 414 552 426 618
rect 1056 552 1068 618
rect 414 546 1068 552
rect 480 518 958 546
rect 480 472 534 518
rect 524 248 534 472
rect 870 472 958 518
rect 870 248 880 472
<< via1 >>
rect 516 2072 1022 2444
rect 1560 1686 1870 1976
rect 72 1136 142 1444
rect 320 1136 390 1444
rect 556 1136 626 1444
rect 792 1136 862 1444
rect 1026 1136 1096 1444
rect 1264 1136 1334 1444
rect 194 766 262 1042
rect 438 768 506 1044
rect 676 768 744 1044
rect 912 774 980 1050
rect 1146 770 1214 1046
rect 426 552 1056 618
rect 534 248 870 518
<< metal2 >>
rect 494 2460 1038 2470
rect 494 2054 1038 2064
rect 520 1970 1020 2054
rect 1560 1976 1870 1986
rect 520 1686 1560 1970
rect 1870 1686 1876 1970
rect 520 1680 1876 1686
rect 520 1482 1020 1680
rect 1560 1676 1870 1680
rect 88 1454 146 1458
rect 326 1454 386 1466
rect 520 1454 1128 1482
rect 72 1444 1338 1454
rect 142 1140 320 1444
rect 72 1126 142 1136
rect 390 1140 556 1444
rect 320 1126 390 1136
rect 626 1140 792 1444
rect 556 1126 626 1136
rect 862 1140 1026 1444
rect 792 1126 862 1136
rect 1096 1140 1264 1444
rect 1026 1126 1096 1136
rect 1334 1140 1338 1444
rect 1264 1126 1334 1136
rect 1264 1124 1322 1126
rect 194 1042 262 1052
rect 438 1044 506 1054
rect 262 768 438 1042
rect 676 1044 744 1054
rect 506 768 676 1042
rect 912 1050 980 1060
rect 744 774 912 1042
rect 1146 1046 1214 1056
rect 980 774 1146 1042
rect 744 770 1146 774
rect 1214 770 1222 1042
rect 744 768 1222 770
rect 262 766 1222 768
rect 194 758 1222 766
rect 194 756 262 758
rect 456 638 956 758
rect 444 628 1008 638
rect 426 618 1056 628
rect 426 542 1056 552
rect 480 518 956 542
rect 480 388 534 518
rect 484 248 534 388
rect 870 248 956 518
rect 484 210 956 248
<< via2 >>
rect 494 2444 1038 2460
rect 494 2072 516 2444
rect 516 2072 1022 2444
rect 1022 2072 1038 2444
rect 494 2064 1038 2072
<< metal3 >>
rect 484 2460 1048 2465
rect 484 2064 494 2460
rect 1038 2064 1048 2460
rect 484 2059 1048 2064
use sky130_fd_pr__nfet_01v8_WUV6BX  XM1
timestamp 1705403419
transform 1 0 704 0 1 1107
box -757 -560 757 560
use sky130_fd_pr__res_xhigh_po_2p85_53STJD  XR2
timestamp 1705403419
transform -1 0 777 0 1 2609
box -451 -725 451 725
<< labels >>
flabel via1 1602 1702 1802 1902 0 FreeSans 256 0 0 0 out
port 0 nsew
flabel metal1 -300 988 -100 1188 0 FreeSans 256 0 0 0 inp
port 1 nsew
flabel metal1 622 3400 822 3600 0 FreeSans 256 180 0 0 vdd
port 2 nsew
flabel via1 620 274 820 474 0 FreeSans 256 0 0 0 vss
port 3 nsew
<< end >>
