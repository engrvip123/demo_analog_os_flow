magic
tech sky130A
magscale 1 2
timestamp 1705403419
<< error_p >>
rect -560 422 -502 428
rect -442 422 -384 428
rect -324 422 -266 428
rect -206 422 -148 428
rect -88 422 -30 428
rect 30 422 88 428
rect 148 422 206 428
rect 266 422 324 428
rect 384 422 442 428
rect 502 422 560 428
rect -560 388 -548 422
rect -442 388 -430 422
rect -324 388 -312 422
rect -206 388 -194 422
rect -88 388 -76 422
rect 30 388 42 422
rect 148 388 160 422
rect 266 388 278 422
rect 384 388 396 422
rect 502 388 514 422
rect -560 382 -502 388
rect -442 382 -384 388
rect -324 382 -266 388
rect -206 382 -148 388
rect -88 382 -30 388
rect 30 382 88 388
rect 148 382 206 388
rect 266 382 324 388
rect 384 382 442 388
rect 502 382 560 388
rect -560 -388 -502 -382
rect -442 -388 -384 -382
rect -324 -388 -266 -382
rect -206 -388 -148 -382
rect -88 -388 -30 -382
rect 30 -388 88 -382
rect 148 -388 206 -382
rect 266 -388 324 -382
rect 384 -388 442 -382
rect 502 -388 560 -382
rect -560 -422 -548 -388
rect -442 -422 -430 -388
rect -324 -422 -312 -388
rect -206 -422 -194 -388
rect -88 -422 -76 -388
rect 30 -422 42 -388
rect 148 -422 160 -388
rect 266 -422 278 -388
rect 384 -422 396 -388
rect 502 -422 514 -388
rect -560 -428 -502 -422
rect -442 -428 -384 -422
rect -324 -428 -266 -422
rect -206 -428 -148 -422
rect -88 -428 -30 -422
rect 30 -428 88 -422
rect 148 -428 206 -422
rect 266 -428 324 -422
rect 384 -428 442 -422
rect 502 -428 560 -422
<< pwell >>
rect -757 -560 757 560
<< nmos >>
rect -561 -350 -501 350
rect -443 -350 -383 350
rect -325 -350 -265 350
rect -207 -350 -147 350
rect -89 -350 -29 350
rect 29 -350 89 350
rect 147 -350 207 350
rect 265 -350 325 350
rect 383 -350 443 350
rect 501 -350 561 350
<< ndiff >>
rect -619 338 -561 350
rect -619 -338 -607 338
rect -573 -338 -561 338
rect -619 -350 -561 -338
rect -501 338 -443 350
rect -501 -338 -489 338
rect -455 -338 -443 338
rect -501 -350 -443 -338
rect -383 338 -325 350
rect -383 -338 -371 338
rect -337 -338 -325 338
rect -383 -350 -325 -338
rect -265 338 -207 350
rect -265 -338 -253 338
rect -219 -338 -207 338
rect -265 -350 -207 -338
rect -147 338 -89 350
rect -147 -338 -135 338
rect -101 -338 -89 338
rect -147 -350 -89 -338
rect -29 338 29 350
rect -29 -338 -17 338
rect 17 -338 29 338
rect -29 -350 29 -338
rect 89 338 147 350
rect 89 -338 101 338
rect 135 -338 147 338
rect 89 -350 147 -338
rect 207 338 265 350
rect 207 -338 219 338
rect 253 -338 265 338
rect 207 -350 265 -338
rect 325 338 383 350
rect 325 -338 337 338
rect 371 -338 383 338
rect 325 -350 383 -338
rect 443 338 501 350
rect 443 -338 455 338
rect 489 -338 501 338
rect 443 -350 501 -338
rect 561 338 619 350
rect 561 -338 573 338
rect 607 -338 619 338
rect 561 -350 619 -338
<< ndiffc >>
rect -607 -338 -573 338
rect -489 -338 -455 338
rect -371 -338 -337 338
rect -253 -338 -219 338
rect -135 -338 -101 338
rect -17 -338 17 338
rect 101 -338 135 338
rect 219 -338 253 338
rect 337 -338 371 338
rect 455 -338 489 338
rect 573 -338 607 338
<< psubdiff >>
rect -721 490 -625 524
rect 625 490 721 524
rect -721 428 -687 490
rect 687 428 721 490
rect -721 -490 -687 -428
rect 687 -490 721 -428
rect -721 -524 -625 -490
rect 625 -524 721 -490
<< psubdiffcont >>
rect -625 490 625 524
rect -721 -428 -687 428
rect 687 -428 721 428
rect -625 -524 625 -490
<< poly >>
rect -564 422 -498 438
rect -564 388 -548 422
rect -514 388 -498 422
rect -564 372 -498 388
rect -446 422 -380 438
rect -446 388 -430 422
rect -396 388 -380 422
rect -446 372 -380 388
rect -328 422 -262 438
rect -328 388 -312 422
rect -278 388 -262 422
rect -328 372 -262 388
rect -210 422 -144 438
rect -210 388 -194 422
rect -160 388 -144 422
rect -210 372 -144 388
rect -92 422 -26 438
rect -92 388 -76 422
rect -42 388 -26 422
rect -92 372 -26 388
rect 26 422 92 438
rect 26 388 42 422
rect 76 388 92 422
rect 26 372 92 388
rect 144 422 210 438
rect 144 388 160 422
rect 194 388 210 422
rect 144 372 210 388
rect 262 422 328 438
rect 262 388 278 422
rect 312 388 328 422
rect 262 372 328 388
rect 380 422 446 438
rect 380 388 396 422
rect 430 388 446 422
rect 380 372 446 388
rect 498 422 564 438
rect 498 388 514 422
rect 548 388 564 422
rect 498 372 564 388
rect -561 350 -501 372
rect -443 350 -383 372
rect -325 350 -265 372
rect -207 350 -147 372
rect -89 350 -29 372
rect 29 350 89 372
rect 147 350 207 372
rect 265 350 325 372
rect 383 350 443 372
rect 501 350 561 372
rect -561 -372 -501 -350
rect -443 -372 -383 -350
rect -325 -372 -265 -350
rect -207 -372 -147 -350
rect -89 -372 -29 -350
rect 29 -372 89 -350
rect 147 -372 207 -350
rect 265 -372 325 -350
rect 383 -372 443 -350
rect 501 -372 561 -350
rect -564 -388 -498 -372
rect -564 -422 -548 -388
rect -514 -422 -498 -388
rect -564 -438 -498 -422
rect -446 -388 -380 -372
rect -446 -422 -430 -388
rect -396 -422 -380 -388
rect -446 -438 -380 -422
rect -328 -388 -262 -372
rect -328 -422 -312 -388
rect -278 -422 -262 -388
rect -328 -438 -262 -422
rect -210 -388 -144 -372
rect -210 -422 -194 -388
rect -160 -422 -144 -388
rect -210 -438 -144 -422
rect -92 -388 -26 -372
rect -92 -422 -76 -388
rect -42 -422 -26 -388
rect -92 -438 -26 -422
rect 26 -388 92 -372
rect 26 -422 42 -388
rect 76 -422 92 -388
rect 26 -438 92 -422
rect 144 -388 210 -372
rect 144 -422 160 -388
rect 194 -422 210 -388
rect 144 -438 210 -422
rect 262 -388 328 -372
rect 262 -422 278 -388
rect 312 -422 328 -388
rect 262 -438 328 -422
rect 380 -388 446 -372
rect 380 -422 396 -388
rect 430 -422 446 -388
rect 380 -438 446 -422
rect 498 -388 564 -372
rect 498 -422 514 -388
rect 548 -422 564 -388
rect 498 -438 564 -422
<< polycont >>
rect -548 388 -514 422
rect -430 388 -396 422
rect -312 388 -278 422
rect -194 388 -160 422
rect -76 388 -42 422
rect 42 388 76 422
rect 160 388 194 422
rect 278 388 312 422
rect 396 388 430 422
rect 514 388 548 422
rect -548 -422 -514 -388
rect -430 -422 -396 -388
rect -312 -422 -278 -388
rect -194 -422 -160 -388
rect -76 -422 -42 -388
rect 42 -422 76 -388
rect 160 -422 194 -388
rect 278 -422 312 -388
rect 396 -422 430 -388
rect 514 -422 548 -388
<< locali >>
rect -721 490 -625 524
rect 625 490 721 524
rect -721 428 -687 490
rect 687 428 721 490
rect -564 388 -548 422
rect -514 388 -498 422
rect -446 388 -430 422
rect -396 388 -380 422
rect -328 388 -312 422
rect -278 388 -262 422
rect -210 388 -194 422
rect -160 388 -144 422
rect -92 388 -76 422
rect -42 388 -26 422
rect 26 388 42 422
rect 76 388 92 422
rect 144 388 160 422
rect 194 388 210 422
rect 262 388 278 422
rect 312 388 328 422
rect 380 388 396 422
rect 430 388 446 422
rect 498 388 514 422
rect 548 388 564 422
rect -607 338 -573 354
rect -607 -354 -573 -338
rect -489 338 -455 354
rect -489 -354 -455 -338
rect -371 338 -337 354
rect -371 -354 -337 -338
rect -253 338 -219 354
rect -253 -354 -219 -338
rect -135 338 -101 354
rect -135 -354 -101 -338
rect -17 338 17 354
rect -17 -354 17 -338
rect 101 338 135 354
rect 101 -354 135 -338
rect 219 338 253 354
rect 219 -354 253 -338
rect 337 338 371 354
rect 337 -354 371 -338
rect 455 338 489 354
rect 455 -354 489 -338
rect 573 338 607 354
rect 573 -354 607 -338
rect -564 -422 -548 -388
rect -514 -422 -498 -388
rect -446 -422 -430 -388
rect -396 -422 -380 -388
rect -328 -422 -312 -388
rect -278 -422 -262 -388
rect -210 -422 -194 -388
rect -160 -422 -144 -388
rect -92 -422 -76 -388
rect -42 -422 -26 -388
rect 26 -422 42 -388
rect 76 -422 92 -388
rect 144 -422 160 -388
rect 194 -422 210 -388
rect 262 -422 278 -388
rect 312 -422 328 -388
rect 380 -422 396 -388
rect 430 -422 446 -388
rect 498 -422 514 -388
rect 548 -422 564 -388
rect -721 -490 -687 -428
rect 687 -490 721 -428
rect -721 -524 -625 -490
rect 625 -524 721 -490
<< viali >>
rect -548 388 -514 422
rect -430 388 -396 422
rect -312 388 -278 422
rect -194 388 -160 422
rect -76 388 -42 422
rect 42 388 76 422
rect 160 388 194 422
rect 278 388 312 422
rect 396 388 430 422
rect 514 388 548 422
rect -607 -338 -573 338
rect -489 -338 -455 338
rect -371 -338 -337 338
rect -253 -338 -219 338
rect -135 -338 -101 338
rect -17 -338 17 338
rect 101 -338 135 338
rect 219 -338 253 338
rect 337 -338 371 338
rect 455 -338 489 338
rect 573 -338 607 338
rect -548 -422 -514 -388
rect -430 -422 -396 -388
rect -312 -422 -278 -388
rect -194 -422 -160 -388
rect -76 -422 -42 -388
rect 42 -422 76 -388
rect 160 -422 194 -388
rect 278 -422 312 -388
rect 396 -422 430 -388
rect 514 -422 548 -388
<< metal1 >>
rect -560 422 -502 428
rect -560 388 -548 422
rect -514 388 -502 422
rect -560 382 -502 388
rect -442 422 -384 428
rect -442 388 -430 422
rect -396 388 -384 422
rect -442 382 -384 388
rect -324 422 -266 428
rect -324 388 -312 422
rect -278 388 -266 422
rect -324 382 -266 388
rect -206 422 -148 428
rect -206 388 -194 422
rect -160 388 -148 422
rect -206 382 -148 388
rect -88 422 -30 428
rect -88 388 -76 422
rect -42 388 -30 422
rect -88 382 -30 388
rect 30 422 88 428
rect 30 388 42 422
rect 76 388 88 422
rect 30 382 88 388
rect 148 422 206 428
rect 148 388 160 422
rect 194 388 206 422
rect 148 382 206 388
rect 266 422 324 428
rect 266 388 278 422
rect 312 388 324 422
rect 266 382 324 388
rect 384 422 442 428
rect 384 388 396 422
rect 430 388 442 422
rect 384 382 442 388
rect 502 422 560 428
rect 502 388 514 422
rect 548 388 560 422
rect 502 382 560 388
rect -613 338 -567 350
rect -613 -338 -607 338
rect -573 -338 -567 338
rect -613 -350 -567 -338
rect -495 338 -449 350
rect -495 -338 -489 338
rect -455 -338 -449 338
rect -495 -350 -449 -338
rect -377 338 -331 350
rect -377 -338 -371 338
rect -337 -338 -331 338
rect -377 -350 -331 -338
rect -259 338 -213 350
rect -259 -338 -253 338
rect -219 -338 -213 338
rect -259 -350 -213 -338
rect -141 338 -95 350
rect -141 -338 -135 338
rect -101 -338 -95 338
rect -141 -350 -95 -338
rect -23 338 23 350
rect -23 -338 -17 338
rect 17 -338 23 338
rect -23 -350 23 -338
rect 95 338 141 350
rect 95 -338 101 338
rect 135 -338 141 338
rect 95 -350 141 -338
rect 213 338 259 350
rect 213 -338 219 338
rect 253 -338 259 338
rect 213 -350 259 -338
rect 331 338 377 350
rect 331 -338 337 338
rect 371 -338 377 338
rect 331 -350 377 -338
rect 449 338 495 350
rect 449 -338 455 338
rect 489 -338 495 338
rect 449 -350 495 -338
rect 567 338 613 350
rect 567 -338 573 338
rect 607 -338 613 338
rect 567 -350 613 -338
rect -560 -388 -502 -382
rect -560 -422 -548 -388
rect -514 -422 -502 -388
rect -560 -428 -502 -422
rect -442 -388 -384 -382
rect -442 -422 -430 -388
rect -396 -422 -384 -388
rect -442 -428 -384 -422
rect -324 -388 -266 -382
rect -324 -422 -312 -388
rect -278 -422 -266 -388
rect -324 -428 -266 -422
rect -206 -388 -148 -382
rect -206 -422 -194 -388
rect -160 -422 -148 -388
rect -206 -428 -148 -422
rect -88 -388 -30 -382
rect -88 -422 -76 -388
rect -42 -422 -30 -388
rect -88 -428 -30 -422
rect 30 -388 88 -382
rect 30 -422 42 -388
rect 76 -422 88 -388
rect 30 -428 88 -422
rect 148 -388 206 -382
rect 148 -422 160 -388
rect 194 -422 206 -388
rect 148 -428 206 -422
rect 266 -388 324 -382
rect 266 -422 278 -388
rect 312 -422 324 -388
rect 266 -428 324 -422
rect 384 -388 442 -382
rect 384 -422 396 -388
rect 430 -422 442 -388
rect 384 -428 442 -422
rect 502 -388 560 -382
rect 502 -422 514 -388
rect 548 -422 560 -388
rect 502 -428 560 -422
<< properties >>
string FIXED_BBOX -704 -507 704 507
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 3.5 l 0.3 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
