magic
tech sky130A
magscale 1 2
timestamp 1705560353
<< locali >>
rect 1072 1600 1156 1886
<< viali >>
rect 450 540 902 618
<< metal1 >>
rect 498 2764 944 3694
rect 464 2002 474 2360
rect 1000 2002 1010 2360
rect -272 1564 248 1566
rect -272 1490 1286 1564
rect -268 1208 -118 1490
rect 118 1486 1286 1490
rect -598 870 -118 1208
rect 64 1088 74 1448
rect 142 1088 152 1448
rect 310 1082 320 1442
rect 388 1082 398 1442
rect 548 1076 558 1436
rect 626 1076 636 1436
rect 782 1076 792 1436
rect 860 1076 870 1436
rect 1018 1078 1028 1438
rect 1096 1078 1106 1438
rect 1252 1078 1262 1438
rect 1330 1078 1340 1438
rect 1524 1142 1534 1414
rect 1770 1142 1780 1414
rect -268 726 -118 870
rect 196 762 206 1010
rect 264 762 274 1010
rect 428 768 438 1016
rect 496 768 506 1016
rect 668 766 678 1014
rect 736 766 746 1014
rect 902 760 912 1008
rect 970 760 980 1008
rect 1132 760 1142 1008
rect 1200 760 1210 1008
rect 248 726 1266 728
rect -272 662 1266 726
rect -272 650 248 662
rect 438 618 914 624
rect 438 540 450 618
rect 902 540 914 618
rect 438 534 914 540
rect 514 516 866 534
rect 514 502 554 516
rect 544 294 554 502
rect 814 502 866 516
rect 814 294 824 502
<< via1 >>
rect 474 2002 1000 2360
rect 74 1088 142 1448
rect 320 1082 388 1442
rect 558 1076 626 1436
rect 792 1076 860 1436
rect 1028 1078 1096 1438
rect 1262 1078 1330 1438
rect 1534 1142 1770 1414
rect 206 762 264 1010
rect 438 768 496 1016
rect 678 766 736 1014
rect 912 760 970 1008
rect 1142 760 1200 1008
rect 450 540 902 618
rect 554 294 814 516
<< metal2 >>
rect 474 2366 1000 2370
rect 422 2360 1024 2366
rect 422 2002 474 2360
rect 1000 2002 1024 2360
rect 422 1480 1024 2002
rect 74 1448 142 1458
rect 422 1456 1092 1480
rect 364 1452 1092 1456
rect 70 1088 74 1430
rect 320 1448 1092 1452
rect 320 1442 1096 1448
rect 142 1088 320 1430
rect 70 1086 320 1088
rect 74 1078 142 1086
rect 388 1438 1096 1442
rect 388 1436 1028 1438
rect 388 1086 558 1436
rect 320 1072 388 1082
rect 626 1086 792 1436
rect 558 1066 626 1076
rect 860 1086 1028 1436
rect 792 1066 860 1076
rect 1262 1438 1330 1448
rect 1096 1086 1262 1430
rect 1028 1068 1096 1078
rect 1534 1414 1784 1430
rect 1770 1142 1784 1414
rect 1534 1086 1784 1142
rect 1262 1068 1330 1078
rect 206 1010 264 1020
rect 194 766 206 982
rect 438 1016 496 1026
rect 264 768 438 982
rect 678 1014 736 1024
rect 496 768 678 982
rect 264 766 678 768
rect 912 1008 970 1018
rect 736 766 912 982
rect 206 752 264 762
rect 438 758 822 766
rect 494 730 822 758
rect 1142 1008 1200 1018
rect 970 766 1142 982
rect 912 750 970 760
rect 1200 766 1210 982
rect 1142 750 1200 760
rect 522 628 822 730
rect 450 618 902 628
rect 450 530 902 540
rect 522 516 822 530
rect 522 294 554 516
rect 814 294 822 516
rect 522 286 822 294
rect 554 284 814 286
use sky130_fd_pr__nfet_01v8_WUV6BX  XM1
timestamp 1705560353
transform -1 0 704 0 1 1107
box -757 -560 757 560
use sky130_fd_pr__res_xhigh_po_2p85_53STJD  XR2
timestamp 1705560353
transform 1 0 743 0 1 2541
box -451 -725 451 725
<< labels >>
flabel via1 578 300 778 500 0 FreeSans 256 0 0 0 vss
port 3 nsew
flabel via1 1564 1192 1764 1392 0 FreeSans 256 0 0 0 out
port 0 nsew
flabel metal1 610 3406 810 3606 0 FreeSans 256 0 0 0 vdd
port 2 nsew
flabel metal1 -520 950 -320 1150 0 FreeSans 256 0 0 0 inp
port 1 nsew
<< end >>
