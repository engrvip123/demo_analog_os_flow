magic
tech sky130A
magscale 1 2
timestamp 1705403069
<< checkpaint >>
rect 148 1460 3570 3204
rect -1260 -766 3570 1460
rect -1260 -2460 1460 -766
<< pwell >>
rect 920 1904 960 1926
<< locali >>
rect 430 1598 816 1940
<< viali >>
rect 498 574 936 622
<< metal1 >>
rect 518 3534 528 3766
rect 746 3534 756 3766
rect 428 2762 438 3168
rect 852 2762 862 3168
rect 402 2040 412 2450
rect 918 2040 928 2450
rect 1772 1682 1782 1924
rect 2008 1682 2018 1924
rect -210 1556 140 1562
rect -210 1488 1286 1556
rect -210 1486 140 1488
rect -210 1328 -116 1486
rect -354 1078 -116 1328
rect 72 1156 82 1410
rect 134 1156 144 1410
rect 312 1154 322 1408
rect 374 1154 384 1408
rect 550 1156 560 1410
rect 612 1156 622 1410
rect 782 1156 792 1410
rect 844 1156 854 1410
rect 1022 1156 1032 1410
rect 1084 1156 1094 1410
rect 1262 1148 1272 1402
rect 1324 1148 1334 1402
rect -210 728 -116 1078
rect 196 802 206 996
rect 260 802 270 996
rect 430 794 440 988
rect 494 794 504 988
rect 664 792 674 986
rect 728 792 738 986
rect 900 786 910 980
rect 964 786 974 980
rect 1140 792 1150 986
rect 1204 792 1214 986
rect -212 726 162 728
rect -212 670 1276 726
rect -212 666 162 670
rect 470 564 480 636
rect 954 564 964 636
rect 588 450 788 458
rect 582 274 592 450
rect 782 274 792 450
rect 588 258 788 274
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
<< via1 >>
rect 528 3534 746 3766
rect 438 2762 852 3168
rect 412 2040 918 2450
rect 1782 1682 2008 1924
rect 82 1156 134 1410
rect 322 1154 374 1408
rect 560 1156 612 1410
rect 792 1156 844 1410
rect 1032 1156 1084 1410
rect 1272 1148 1324 1402
rect 206 802 260 996
rect 440 794 494 988
rect 674 792 728 986
rect 910 786 964 980
rect 1150 792 1204 986
rect 480 622 954 636
rect 480 574 498 622
rect 498 574 936 622
rect 936 574 954 622
rect 480 564 954 574
rect 592 274 782 450
<< metal2 >>
rect 400 3832 896 3858
rect 392 3766 896 3832
rect 392 3534 528 3766
rect 746 3534 896 3766
rect 392 3168 896 3534
rect 392 2766 438 3168
rect 400 2762 438 2766
rect 852 2762 896 3168
rect 400 2752 896 2762
rect 412 2456 918 2460
rect 408 2450 922 2456
rect 408 2040 412 2450
rect 918 2040 922 2450
rect 408 1926 922 2040
rect 1782 1926 2008 1934
rect 408 1924 2034 1926
rect 408 1682 1782 1924
rect 2008 1682 2034 1924
rect 408 1650 2034 1682
rect 82 1410 134 1420
rect 78 1246 82 1408
rect 322 1408 374 1418
rect 408 1410 922 1650
rect 408 1408 560 1410
rect 134 1246 322 1408
rect 82 1146 134 1156
rect 374 1246 560 1408
rect 322 1144 374 1154
rect 612 1246 792 1410
rect 560 1146 612 1156
rect 844 1408 922 1410
rect 1032 1410 1084 1420
rect 844 1246 1032 1408
rect 792 1146 844 1156
rect 1272 1408 1324 1412
rect 1084 1402 1330 1408
rect 1084 1246 1272 1402
rect 1032 1146 1084 1156
rect 1324 1246 1330 1402
rect 1272 1138 1324 1148
rect 206 996 260 1006
rect 198 802 206 978
rect 440 988 494 998
rect 260 802 440 978
rect 198 798 440 802
rect 206 792 260 798
rect 674 986 728 996
rect 494 798 674 978
rect 440 784 494 794
rect 558 792 674 798
rect 910 980 964 990
rect 728 798 910 978
rect 728 792 878 798
rect 558 646 878 792
rect 1150 986 1204 996
rect 964 798 1150 978
rect 910 776 964 786
rect 1204 798 1208 978
rect 1150 782 1204 792
rect 480 636 954 646
rect 480 554 954 564
rect 558 450 878 554
rect 558 274 592 450
rect 782 274 878 450
rect 558 262 878 274
use sky130_fd_pr__res_xhigh_po_2p85_RYTYPJ  sky130_fd_pr__res_xhigh_po_2p85_RYTYPJ_0
timestamp 1695730206
transform -1 0 659 0 1 2613
box -451 -741 451 741
use sky130_fd_pr__nfet_01v8_WUV6BX  XM1
timestamp 1695627866
transform 1 0 704 0 1 1107
box -757 -560 757 560
use sky130_fd_pr__res_xhigh_po_2p85_53STJD  XR2
timestamp 0
transform 1 0 1859 0 1 1219
box -451 -725 451 725
<< labels >>
flabel via1 1800 1710 2000 1910 0 FreeSans 256 0 0 0 out
port 1 nsew
flabel metal1 588 258 788 458 0 FreeSans 256 0 0 0 vss
port 3 nsew
flabel metal1 -342 1102 -142 1302 0 FreeSans 256 0 0 0 inp
port 0 nsew
flabel via1 540 3546 740 3746 0 FreeSans 256 0 0 0 vdd
port 2 nsew
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 out
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 inp
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 vdd
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 vss
<< end >>
