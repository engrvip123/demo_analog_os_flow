magic
tech sky130A
magscale 1 2
timestamp 1705560353
<< pwell >>
rect -451 -725 451 725
<< psubdiff >>
rect -415 655 -319 689
rect 319 655 415 689
rect -415 593 -381 655
rect 381 593 415 655
rect -415 -655 -381 -593
rect 381 -655 415 -593
rect -415 -689 -319 -655
rect 319 -689 415 -655
<< psubdiffcont >>
rect -319 655 319 689
rect -415 -593 -381 593
rect 381 -593 415 593
rect -319 -689 319 -655
<< xpolycontact >>
rect -285 127 285 559
rect -285 -559 285 -127
<< xpolyres >>
rect -285 -127 285 127
<< locali >>
rect -415 655 -319 689
rect 319 655 415 689
rect -415 593 -381 655
rect 381 593 415 655
rect -415 -655 -381 -593
rect 381 -655 415 -593
rect -415 -689 -319 -655
rect 319 -689 415 -655
<< viali >>
rect -269 144 269 541
rect -269 -541 269 -144
<< metal1 >>
rect -281 541 281 547
rect -281 144 -269 541
rect 269 144 281 541
rect -281 138 281 144
rect -281 -144 281 -138
rect -281 -541 -269 -144
rect 269 -541 281 -144
rect -281 -547 281 -541
<< properties >>
string FIXED_BBOX -398 -672 398 672
string gencell sky130_fd_pr__res_xhigh_po_2p85
string library sky130
string parameters w 2.850 l 1.43 m 1 nx 1 wmin 2.850 lmin 0.50 rho 2000 val 1.135k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 2.850 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
